* Simple opamp, 0.18u, 1.8V, HSPICE

* Any include or lib that is set from PyOPUS (specified in problem definition) 
* must not be specified here. 

* Include files - fixed
.include 'mosmm.inc'

* Any parameter that is set from PyOPUS (specified in problem definition) 
* must not be specified here. 

* Operating conditions - fixed
.param lev1=0
.param lev2=0.5
.param tstart=1e-9
.param tr=1e-9
.param tf=1e-9
.param pw=500e-9
.param ibias=1.000000000000e-004 
.param rfb=1e6
.param rin=1e6

* Design parameters - fixed
.param out_w=4.800592541419e-005
.param out_l=3.750131780858e-007
.param load_w=3.486243671853e-005
.param load_l=2.572996921261e-006
.param dif_w=7.728734451428e-006
.param dif_l=1.082371380389e-006
.param c_out=8.211596855053e-012
.param r_out=1.968986740568e+001

* inp inn out vdd vss bias slp slpx
.subckt amp 3 4 5 1 2 7 11 12
xmp1 9 10 1 1  submodp w=load_w l=load_l m=2
xmp2 10 10 1 1 submodp w=load_w l=load_l m=2
xmp1s 9 12 1 1 submodp w=1u        l=0.5u
xmp3 5 9 1 1   submodp w=out_w   l=out_l   m=16
xmn2 9 3 8 2   submodn w=dif_w   l=dif_l 
xmn3 10 4 8 2  submodn w=dif_w   l=dif_l 
xmn1s 7 11 2 2 submodn w=1u        l=0.5u
xmn1b 7 7 2 2  submodn w=mirr_w  l=mirr_l  m=2
xmn1 8 7 2 2   submodn w=mirr_w  l=mirr_l  m=2
xmn4 5 7 2 2   submodn w=mirr_w  l=mirr_l  m=16
cout 5a 9 c=c_out
rout 5 5a r=r_out
.ends

* Test topology
x1 inp inn out vdd 0 bias 0 vdd amp
vdd vdd 0 dc=vdd
ibias vdd bias dc=ibias
rfb out inn rfb
rin in inn rin
vcom inp 0 dc='vdd/2'
vin in inp dc=0 ac=1 pulse (lev1 lev2 tstart tr tf pw)
rload out 0 100k
cload out 0 0.5p

* This file is included in the main simulator input file. 
* Do not add .end - it is added by PyOPUS to the main input file. 
